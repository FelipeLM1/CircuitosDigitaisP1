-- SUBTRATOR
-- 
--	PEGA OS VALORES INVERTE E SOMA. 
--

